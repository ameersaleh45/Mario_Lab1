library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pic_pipe is
port(
	  ADDR    : in integer range 0 to 4095;
	  Q       : out std_logic_vector(7 downto 0)
);
end pic_pipe;

architecture arch of pic_pipe is

type matrix is array(0 to 4095) of std_logic_vector(7 downto 0);

constant pipe : matrix := (
							X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
							X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"00", X"00", 
							X"00", X"00", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", 
							X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
							X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13", 
							X"13", X"13", X"13", X"13", X"00", X"00", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"14", X"BC", X"BC", X"14", X"14", X"BC", X"BC", X"BC", X"BC", X"00", X"00", X"13", X"13", X"13", X"13"  
						  );
begin

	Q <= pipe(ADDR);		
			
end arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pic_game_over is
port(
	  ADDR    : in integer range 0 to 4479;
	  Q       : out std_logic_vector(7 downto 0)
);
end pic_game_over;

architecture arch of pic_game_over is

type matrix is array(0 to 4479) of std_logic_vector(7 downto 0);

constant game_over : matrix := (  
X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"FF", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"B6", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"B6", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"B6", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"B6", X"92", X"B6", X"FF", X"FF", X"FF", X"FF", X"DB", X"6D", X"FF", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"FF", X"FF", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"92", X"B6", X"92", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"DB", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"24", X"00", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"6D", X"00", X"6D", X"DB", X"B6", X"B6", X"B6", X"DB", X"B6", X"00", X"00", X"00", X"00", X"DB", X"B6", X"B6", X"B6", X"B6", X"DB", X"24", X"00", X"92", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"B6", X"00", X"00", X"92", X"B6", X"6D", X"DB", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"92", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"DB", X"00", X"00", X"DB", X"B6", X"B6", X"DB", X"00", X"00", X"92", X"DB", X"B6", X"DB", X"6D", X"00", X"6D", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"00", X"24", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"DB", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"DB", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"49", X"49", X"49", X"49", X"49", X"49", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"6D", X"24", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"49", X"49", X"49", X"49", X"49", X"49", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"B6", X"24", X"6D", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"B6", X"24", X"49", X"49", X"49", X"49", X"49", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"24", X"49", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"B6", X"B6", X"DB", X"24", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"DB", X"B6", X"B6", X"B6", X"B6", X"DB", X"B6", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"DB", X"B6", X"B6", X"B6", X"B6", X"B6", X"DB", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"B6", X"49", X"49", X"49", X"49", X"49", X"49", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"B6", X"49", X"49", X"49", X"49", X"49", X"6D", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"DB", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"92", X"6D", X"DB", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"24", X"92", X"92", X"92", X"92", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"00", X"92", X"92", X"92", X"92", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"B6", X"92", X"DB", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"DB", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"6D", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"6D", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"6D", X"6D", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"B6", X"49", X"92", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"B6", X"49", X"92", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"92", X"FF", X"FF", X"FF", X"DB", X"49", X"6D", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"92", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"B6", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"49", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"B6", X"FF", X"FF", X"FF", X"92", X"00", X"6D", X"FF", X"FF", X"FF", X"DB", X"00", X"24", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"00", X"00", X"00", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"00", X"49", X"FF", X"FF", X"FF", X"FF", X"00", X"00", X"FF", X"FF", X"FF", X"FF", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"24", X"B6", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"B6", X"24", X"00", X"B6", X"92", X"92", X"B6", X"00", X"00", X"6D", X"B6", X"92", X"B6", X"6D", X"00", X"49", X"B6", X"92", X"B6", X"6D", X"00", X"24", X"B6", X"92", X"92", X"B6", X"00", X"00", X"B6", X"92", X"92", X"B6", X"24", X"00", X"6D", X"B6", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"00", X"00", X"92", X"B6", X"6D", X"FF", X"FF", X"FF", X"FF", X"92", X"92", X"FF", X"00", X"00", X"6D", X"B6", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"B6", X"00", X"00", X"B6", X"92", X"92", X"92", X"92", X"B6", X"24", X"00", X"00", X"00", X"00", X"00", X"6D", X"B6", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"92", X"B6", X"00", X"24", X"B6", X"92", X"92", X"92", X"00", X"00", X"92", X"92", X"92", X"B6", X"24", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"FF", X"24", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"92", X"B6", X"6D", X"DB", X"FF", X"FF", X"FF", X"92", X"92", X"DB", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"24", X"FF", X"DB", X"FF", 
X"FF", X"DB", X"DB", X"6D", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"DB", X"92", X"92", X"FF", X"FF", X"FF", X"FF", X"92", X"6D", X"FF", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"24", X"FF", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"6D", X"DB", X"DB", X"FF", 
X"FF", X"FF", X"92", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"6D", X"92", X"FF", X"FF", X"FF", X"FF", X"B6", X"6D", X"92", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"92", X"FF", X"FF", 
X"FF", X"FF", X"DB", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"DB", X"FF", X"FF", X"FF", X"FF", X"DB", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"DB", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"B6", X"92", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"92", X"B6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"92", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"92", X"92", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"6D", X"92", X"B6", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"FF", X"FF", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"DB", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF"
 );
begin

	Q <= game_over(ADDR);		
			
end arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pic_ground is
port(
	  ADDR    : in std_logic_vector(11 downto 0);
	  Q       : out std_logic_vector(7 downto 0)
);
end pic_ground;

architecture arch of pic_ground is

type matrix is array(0 to 4095) of std_logic_vector(7 downto 0);

constant ground : matrix := (
X"A8", X"A8", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"05", X"05", X"A9", X"A9", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"A9", X"A8", X"A8", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"05", X"05", X"A9", X"A9", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"93", X"A9", X"A9", X"A8", 
X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", 
X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"F6", 
X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", 
X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", 
X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", 
X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"C8", X"C8", X"C8", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"00", 
X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6", 
X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"00", X"00", X"F6", X"F6", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00", X"00", X"F6"			
							  );
begin

	Q <= ground(to_integer(unsigned(ADDR)));		
			
end arch;
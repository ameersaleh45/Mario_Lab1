library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_arith.all; --

-------------------------------------------------
-- This module contains the static objects of the game, cloubds, blocks, pipes
-- it uses generic object generator and duplicate objects on the screen reading from 
-- a single ROM, uses arrays of coordinates that can be changed easily to create
-- new game levels. it's also scalable, you can add new objects to the game using the
-- generic component
-------------------------------------------------

entity static_objects is
	port 	(
	   	CLK  			: in std_logic; 
		RESETn			: in std_logic;
		
		oCoord_X		: in integer;						 -- current pixel that the VGA controller is handling
		oCoord_Y		: in integer;
		map_offset		: in integer;						 -- current screen game offset from beginning 
		game_over		: in std_logic;						 -- turns on the game_over sign
		start			: in std_logic;						 -- turns on the start sign
		win				: in std_logic;
		show_map		: in std_logic;
		drawing_request					: out std_logic ;					 -- whether an object exists in current pixel
		mVGA_RGB 						: out std_logic_vector(7 downto 0)   -- color of current character pixel in 8bit

	);
	
end static_objects;

architecture behav of static_objects is 

	--------------------------------------------------
	-- roms of the game static objects
	--------------------------------------------------
	
	COMPONENT generic_object IS
		port (
					CLK  			: in std_logic; 
					RESETn			: in std_logic;
					
					oCoord_X		: in integer;						 
					oCoord_Y		: in integer;
					map_offset		: in integer;
					
					ObjectStartX	: in integer;						
					ObjectStartY 	: in integer;
					object_X_size	: in integer;
					object_Y_size 	: in integer;
					
					drawing_request	: out std_logic ;
					address 		: out integer  			
			);
	
	END COMPONENT;
	
	---------------------objects---------------------
	
	constant StartSizeX : integer := 72;
	constant StartSizeY : integer := 35;
	
	COMPONENT pic_start IS
		port(
				ADDR    : in integer range 0 to (StartSizeX*StartSizeY - 1);
				Q       : out std_logic_vector(7 downto 0)
		);
	END COMPONENT;
	
	signal muxed_start				: integer range 0 to (StartSizeX*StartSizeY - 1) := 0;
	signal start_rgb				: std_logic_vector (7 downto 0);
	signal drawing_request_start	: std_logic := '0';
	
	-------------------------------------------------- 
	
	constant winSizeX 		: integer := 82;
	constant winSizeY 		: integer := 35;
	
	COMPONENT pic_win IS
		port(
			ADDR    : in integer range 0 to (winSizeX*winSizeY - 1);
			Q       : out std_logic_vector(7 downto 0)
		);
	END COMPONENT;
	
	signal muxed_win					: integer range 0 to (winSizeX*winSizeY - 1) := 0;
	signal win_rgb						: std_logic_vector (7 downto 0);
	signal drawing_request_win			: std_logic := '0';	
	-------------------------------------------------- 
	
	constant GameOverSizeX 		: integer := 128;
	constant GameOverSizeY 		: integer := 35;
	
	COMPONENT pic_game_over IS
		port(
			ADDR    : in integer range 0 to (GameOverSizeX*GameOverSizeY - 1);
			Q       : out std_logic_vector(7 downto 0)
		);
	END COMPONENT;
	
	signal muxed_game_over				: integer range 0 to (GameOverSizeX*GameOverSizeY - 1) := 0;
	signal game_over_rgb				: std_logic_vector (7 downto 0);
	signal drawing_request_game_over	: std_logic := '0';
	
	-------------------------------------------------- 
	
	constant CastleSizeX : integer := 54;
	constant CastleSizeY : integer := 64;
	
	COMPONENT pic_castle IS
		port(
			  ADDR    : in integer range 0 to (CastleSizeX*CastleSizeY - 1);
			  Q       : out std_logic_vector(7 downto 0)
		);
	END COMPONENT;
	
	signal muxed_castle				: integer range 0 to (CastleSizeX*CastleSizeY - 1) := 0;
	signal castle_rgb	 			: std_logic_vector (7 downto 0);
	signal drawing_request_castle	: std_logic := '0';
	
	-------------------------------------------------- 
	
	constant bigCloudSizeX : integer := 96;
	constant bigCloudSizeY : integer := 48;
	
	COMPONENT pic_big_cloud IS
		PORT
		(
		    ADDR    	: in integer range 0 to (bigCloudSizeX*bigCloudSizeY - 1);
			q			: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
	END COMPONENT;
	
	
	signal muxed_big_cloud 			: integer range 0 to (bigCloudSizeX*bigCloudSizeY - 1) := 0;
	signal big_cloud_rgb  			: std_logic_vector (7 downto 0);	
	signal drawing_request_bCloud	: std_logic := '0';
	
	-------------------------------------------------- 	
	
	constant smallCloudSizeX : integer := 64;
	constant smallCloudSizeY : integer := 48;
	
	COMPONENT pic_small_cloud IS
		PORT
		(
		    ADDR    	: in integer range 0 to (smallCloudSizeX*smallCloudSizeY - 1);
			q			: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
	END COMPONENT;
	
	
	signal muxed_small_cloud		: integer range 0 to (smallCloudSizeX*smallCloudSizeY - 1) := 0;
	signal small_cloud_rgb 	 		: std_logic_vector (7 downto 0);
	signal drawing_request_sCloud	: std_logic := '0';
	
	-------------------------------------------------- 	
	
	constant brickSizeX : integer := 32;
	constant brickSizeY : integer := 32;
	
	COMPONENT pic_brick IS
		PORT
		(
		    ADDR    	: in integer range 0 to (brickSizeX*brickSizeY - 1);
			q			: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
	END COMPONENT;
		
	signal muxed_brick 				: integer range 0 to (brickSizeX*brickSizeY - 1) := 0;
	signal brick_rgb 				: std_logic_vector (7 downto 0);
	signal drawing_request_brick	: std_logic := '0';
	
	-------------------------------------------------- 	
	
	constant pipeSizeX : integer := 64;
	constant pipeSizeY : integer := 64;
	
	COMPONENT pic_pipe IS
		PORT
		(
		    ADDR    	: in integer range 0 to (pipeSizeX*pipeSizeY - 1);
			q			: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
	END COMPONENT;	
	
	signal muxed_pipe  				: integer range 0 to (pipeSizeX*pipeSizeY - 1) := 0;
	signal pipe_rgb	   				: std_logic_vector (7 downto 0);
	signal drawing_request_pipe		: std_logic := '0';
	
	--------------------------------------------------
	-- creating a map
	--------------------------------------------------
	
	signal drawing_request_sig	: std_logic := '0';				-- global drawing request
	
	type drawing_requests_array			 is array (0 to 9) of std_logic;
	type addresses_array				 is array (0 to 9) of integer;
	
	type drawing_requests_array9		 is array (1 to 9) of std_logic;
	type addresses_array9				 is array (1 to 9) of integer;

	signal address_start 				 : integer := 0;
	signal address_game_over 			 : integer := 0;
	signal address_castle 				 : integer := 0;
	signal address_win 					 : integer := 0;

	-----------------------------------------------------
	-- arrays containing coordinates 
	-----------------------------------------------------
	type object_locations			 is array (0 to 9) of integer;
	type object_locations9			 is array (1 to 9) of integer;
	constant H0					: integer := 416;
	constant H1					: integer := 288;
	constant H2					: integer := 145;

	
	--------------------------------------------------------------------------------------------------------
	constant small_clouds_locsX			: object_locations 			:= (50, 300,3000 ,680,3500,1100,1300,1650,2150,2600);
	constant small_clouds_locsY			: object_locations 			:= (18, 23, 22 , 22, 25, 23, 25 ,64, 50, 56 );
	signal small_clouds_addresses		: addresses_array 			:= ( others => 0 );
	signal small_clouds_dr	 			: drawing_requests_array 	:= ( others => '0' );
	
	--------------------------------------------------------------------------------------------------------
	constant big_clouds_locsX	 		: object_locations 			:= (150,1820,2000,1000, 1200,1450,2300,2800,3900,3600 );
	constant big_clouds_locsY	 		: object_locations 			:= ( 52,52,52,52,52,52,52,52,52,52);
	signal big_clouds_addresses			: addresses_array 			:= ( others => 0 );
	signal big_clouds_dr	 			: drawing_requests_array 	:= ( others => '0' );
	
	--------------------------------------------------------------------------------------------------------
	constant bricks_locsX1	 			: object_locations 			:= (24,28,32,50,54,77,81,96,100,146);
	constant bricks_locsY1	 			: object_locations 			:= (9,9,9,7,7,9,9,7,7,9);
	constant bricks_locsX2	 			: object_locations 			:= (150,190,194,220,230,260,324,304,308,320);
	constant bricks_locsY2	 			: object_locations 			:= (9,9,9,9,7,9,9,7,7,9);
	signal bricks_addresses1 			: addresses_array 			:= ( others => 0 );
	signal bricks_dr1 		 			: drawing_requests_array 	:= ( others => '0' );
	signal bricks_addresses2 			: addresses_array 			:= ( others => 0 );
	signal bricks_dr2 		 			: drawing_requests_array 	:= ( others => '0' );
	
	--------------------------------------------------------------------------------------------------------
	constant pipes_locsX				: object_locations 			:= (124,168,200,300,350,350,350,350,350,350);
	constant pipes_locsY				: object_locations 			:= (11,11,11,11,11,11,11,11,11,11);	
	signal pipes_addresses				: addresses_array  			:= ( others => 0 );
	signal pipes_dr 		 			: drawing_requests_array 	:= ( others => '0' );
	
	--------------------------------------------------------------------------------------------------------
	constant CrazyBricks_locsX	 		: object_locations9 		:= (1,6,12 ,          0,7,11,      1,7,11);
	constant CrazyBricks_locsY	 		: object_locations9 		:= (H0,H0,H0 ,        H1,H1,H1,    H2,H2,H2);
	signal crazy_bricks_addresses		: addresses_array9 			:= ( others => 0 );
	signal crazyBricks_dr 	 			: drawing_requests_array9 	:= ( others => '0' );
	
	
	signal CblockAppear					: std_logic_vector(9 downto 1) := (others => '1' );
	
	-- objects are placed in coordinates that are a multiplier of the moving speed so the collisions would be identified immediately
	constant objectXMultiplier : integer := 8;	
	constant objectYMultiplier  : integer := 32;
	constant crazybrickMultiplier: integer := 32;
	constant crazy_level_offset : integer := 3000;
	
	-----------------------------------------------------
	--------------------------------------------------------------------------------------------------------
	----------------------------------------MOST AWESOME FEATURE YET----------------------------------------
	--------------------------------------------------------------------------------------------------------
	
	type matrix is array(0 to 4127) of std_logic_vector(7 downto 0);
	signal small_map : matrix := ( 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00",
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"00", 
X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00",
X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00",
X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00",
X"00", X"00", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"C8", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"	
	); 
	
	signal first_cycle : std_logic := '1'; -- indicates first cycle of the game, we want to create the small map once
	constant mapSizeX 			: integer := 129;
	constant mapSizeY 			: integer := 32;
	signal address_map 		    : integer := 0;
	signal drawing_request_map	: std_logic := '0';
	--------------------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------------------
	
	
	component random_ctr3   is
	port (
		CLK 		: in 	std_logic;
		RESETN 		: in 	std_logic; 
		
        random1	 	: out 	std_logic_vector (2 downto 0);
        random2	 	: out 	std_logic_vector (2 downto 0);
        random3	 	: out 	std_logic_vector (2 downto 0) 

    );
	end component;
	
	signal rand1 : std_logic_vector (2 downto 0);
	signal rand2 : std_logic_vector (2 downto 0);
	signal rand3 : std_logic_vector (2 downto 0);
	
	component dividerT is	--one HZ clk
	port (
		CLK 		: in 	std_logic; --Clock, active high
        RESETN 		: in 	std_logic; --Async. Reset, active low
        HZ			: in 	integer;
        speed		: in    integer;
        rate		: in 	integer;
        slowClk 	: out 	std_logic -- output CLK
    );
	end component;
	constant Hz 	 : integer := 51234567;
	signal HZclk : std_logic;
	-----------------------------------------------------

	
	begin
		
		-- one rom per object, multiple readers
				
		small_cloud_rom  	: pic_small_cloud 		port map(muxed_small_cloud,small_cloud_rgb);
		big_cloud_rom		: pic_big_cloud			port map(muxed_big_cloud,big_cloud_rgb);
		brick_rom			: pic_brick				port map(muxed_brick,brick_rgb);
		pipe_rom			: pic_pipe  			port map(muxed_pipe,pipe_rgb);
		start_rom			: pic_start				port map(muxed_start,start_rgb);
		game_over_rom		: pic_game_over			port map(muxed_game_over,game_over_rgb);
		castle_rom			: pic_castle			port map(muxed_castle,castle_rgb);
		win_rom				: pic_win				port map(muxed_win,win_rgb);
		
		-----------------------------------------------------------------
		-- static objects of the game --TODO make semi-random generations
		-----------------------------------------------------------------
		HZclk1 		: dividerT 		 port map(CLK, RESETn, Hz ,0,0, HZclk);
		random		: random_ctr3 	 port map(CLK, RESETn,rand1,rand2,rand3);
		
		start1		: generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,282, 180, StartSizeX,  StartSizeY,drawing_request_start, address_start);
		game_over1	: generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,256+map_offset, 180, GameOverSizeX, GameOverSizeY ,drawing_request_game_over, address_game_over);
		castle1		: generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,4058 , 353, CastleSizeX, CastleSizeY, drawing_request_castle,address_castle);
		win1		: generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,285+map_offset, 180, winSizeX, winSizeY,drawing_request_win, address_win);
		small_map1	: generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,500+map_offset, 100, mapSizeX, mapSizeY,drawing_request_map, address_map);
		
		small_clouds :		for i in 0 to 9 generate
								small_clouds :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset, small_clouds_locsX(i)  , small_clouds_locsY(i), smallCloudSizeX, smallCloudSizeY, small_clouds_dr(i), small_clouds_addresses(i));
							end generate small_clouds;
		
		
		big_clouds :		for i in 0 to 9 generate
								big_clouds :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset, big_clouds_locsX(i)  , big_clouds_locsY(i), bigCloudSizeX, bigCloudSizeY,big_clouds_dr(i), big_clouds_addresses(i));
							end generate big_clouds;
							
							
		bricks1 :			for i in 0 to 9 generate
								bricks1 :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset, bricks_locsX1(i) * objectXMultiplier  ,  bricks_locsY1(i) * objectYMultiplier , brickSizeX, brickSizeY,bricks_dr1(i), bricks_addresses1(i));
							end generate bricks1;
		
		bricks2 :			for i in 0 to 9 generate
								bricks2 :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset, bricks_locsX2(i) * objectXMultiplier  ,  bricks_locsY2(i) * objectYMultiplier , brickSizeX, brickSizeY,bricks_dr2(i), bricks_addresses2(i));
							end generate bricks2;
		
		pipes :				for i in 0 to 9 generate	
								pipes :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,	pipes_locsX(i) * objectXMultiplier, pipes_locsY(i) * objectYMultiplier, pipeSizeX, pipeSizeY,pipes_dr(i), pipes_addresses(i));
							end generate pipes;
		
		
		crazyLevel :		for i in 1 to 9 generate	
								crazyLevel :generic_object port map(CLK, RESETn, oCoord_X, oCoord_Y, map_offset,CrazyBricks_locsX(i)*crazybrickMultiplier + crazy_level_offset, CrazyBricks_locsY(i), brickSizeX, brickSizeY,crazyBricks_dr(i), crazy_bricks_addresses(i));
							end generate crazyLevel;
		
		
														
		 process ( RESETn, CLK)
			
		   begin
				if RESETn = '0' then
					drawing_request			<= '0' ;				
					mVGA_RGB				<= (others => '0');	
					muxed_small_cloud 		<= 0;
					muxed_big_cloud 		<= 0;
					muxed_brick 			<= 0;
					muxed_pipe 				<= 0;
					muxed_start				<= 0;
					muxed_game_over			<= 0;
					muxed_castle			<= 0;
					muxed_win				<= 0;
					first_cycle 			<= '1';
					
				elsif rising_edge(CLK) then
				
					drawing_request_sig <= '0';
					if(drawing_request_map = '1' and show_map = '1' )then
							drawing_request_sig <= '1';
							mVGA_RGB <= small_map(address_map);		
					elsif(drawing_request_start = '1' and start = '0') then 
							drawing_request_sig <= '1';
							muxed_start <= address_start;
							mVGA_RGB <= start_rgb;				
					elsif(drawing_request_game_over = '1' and game_over = '1') then 
							drawing_request_sig <= '1';
							muxed_game_over <= address_game_over;
							mVGA_RGB <= game_over_rgb;
					elsif(drawing_request_win = '1' and win = '1') then 
							drawing_request_sig <= '1';
							muxed_win <= address_win;
							mVGA_RGB <= win_rgb;
					elsif(drawing_request_castle = '1') then 
							drawing_request_sig <= '1';
							muxed_castle <= address_castle;
							mVGA_RGB <= castle_rgb;
					else
						
						for i in 0 to 9 loop
							if(small_clouds_dr(i) = '1') then 
								drawing_request_sig <= '1';
								muxed_small_cloud <= small_clouds_addresses(i);
								mVGA_RGB <= small_cloud_rgb;
								exit;	
											
							elsif(big_clouds_dr(i) = '1') then 
								drawing_request_sig <= '1';
								muxed_big_cloud <= big_clouds_addresses(i);
								mVGA_RGB <= big_cloud_rgb;
								exit;
								
							elsif(bricks_dr1(i) = '1') then 
								drawing_request_sig <= '1';
								muxed_brick <= bricks_addresses1(i);
								mVGA_RGB <= brick_rgb;
								exit;
									
							elsif(bricks_dr2(i) = '1') then 
								drawing_request_sig <= '1';
								muxed_brick <= bricks_addresses2(i);
								mVGA_RGB <= brick_rgb;
								exit;
								
							elsif(pipes_dr(i) = '1') then 
								drawing_request_sig <= '1';
								muxed_pipe <= pipes_addresses(i);
								mVGA_RGB <= pipe_rgb;
								exit;							
							end if;

						end loop;	
							
						if(HZclk = '1') then
							CblockAppear(9 downto 7)  	<= rand1(2 downto 0);
							CblockAppear(6 downto 4) 	<= rand2(2 downto 0);
							CblockAppear(3 downto 1) 	<= rand3(2 downto 0);
						end if;
						
						for j in 1 to 9 loop
							if(crazyBricks_dr(j) = '1' and CblockAppear(j) = '1') then 
								drawing_request_sig <= '1';
								muxed_brick <= crazy_bricks_addresses(j);
								mVGA_RGB <= brick_rgb; 
								exit;
							end if;				
						end loop;
						
					end if;
					
					drawing_request <= drawing_request_sig;
					
					if(first_cycle = '1') then						
						for i in 0 to 9 loop
							-- bricks
							small_map(129* bricks_locsY1(i)*2 +(bricks_locsX1(i)/4+1)) <= "11001000";
							small_map(129* bricks_locsY2(i)*2 +(bricks_locsX2(i)/4+1)) <= "11001000";
							-- pipes
							small_map(129* pipes_locsY(i)*2 +(pipes_locsX(i)/4+1)) <= "10111100";
							small_map(129* pipes_locsY(i)*2 +(pipes_locsX(i)/4+2)) <= "10111100";
							small_map(129* (pipes_locsY(i)+1)*2 +(pipes_locsX(i)/4+1)) <= "10111100";
							small_map(129* (pipes_locsY(i)+1)*2 +(pipes_locsX(i)/4+2)) <= "10111100";
							--small clouds
							small_map(129* (small_clouds_locsY(i)+1)/16 +(small_clouds_locsX(i)/32+1)) <= "11111111";
							small_map(129* (small_clouds_locsY(i)+1)/16 +(small_clouds_locsX(i)/32+2)) <= "11111111";
							small_map(129* ((small_clouds_locsY(i)+1)/16+1) +(small_clouds_locsX(i)/32+1)) <= "11111111";
							small_map(129* ((small_clouds_locsY(i)+1)/16+1)+(small_clouds_locsX(i)/32+2)) <= "11111111";
							--big_clouds
							small_map(129* (big_clouds_locsY(i)+1)/16 +(big_clouds_locsX(i)/32+1)) <= "11111111";
							small_map(129* (big_clouds_locsY(i)+1)/16 +(big_clouds_locsX(i)/32+2)) <= "11111111";
							small_map(129* (big_clouds_locsY(i)+1)/16 +(big_clouds_locsX(i)/32+3)) <= "11111111";
							small_map(129* ((big_clouds_locsY(i)+1)/16+1) +(big_clouds_locsX(i)/32+1)) <= "11111111";
							small_map(129* ((big_clouds_locsY(i)+1)/16+1)+(big_clouds_locsX(i)/32+2)) <= "11111111";
							small_map(129* ((big_clouds_locsY(i)+1)/16+1)+(big_clouds_locsX(i)/32+3)) <= "11111111";
						end loop;
						first_cycle <= '0';
					end if;
				end if;
		 end process;

				
end behav;		
		
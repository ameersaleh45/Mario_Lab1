library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pic_castle is
port(
	  ADDR    : in integer range 0 to 3455;
	  Q       : out std_logic_vector(7 downto 0)
);
end pic_castle;

architecture arch of pic_castle is

type matrix is array(0 to 3455) of std_logic_vector(7 downto 0);

constant castle : matrix := (
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"D1", X"F6", X"13", X"13", X"13", X"CD", X"CD", X"13", X"13", X"13", X"D1", X"CD", X"CD", X"13", X"13", X"13", X"CD", X"D6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"C8", X"F1", X"13", X"13", X"13", X"C4", X"C4", X"13", X"13", X"13", X"CC", X"C4", X"C8", X"13", X"13", X"13", X"C4", X"D1", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"68", X"D2", X"13", X"13", X"13", X"40", X"40", X"13", X"13", X"13", X"88", X"40", X"64", X"13", X"13", X"13", X"40", X"8D", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"ED", X"C8", X"A4", X"80", X"E8", X"A4", X"C8", X"E8", X"60", X"A4", X"E8", X"64", X"E8", X"E8", X"40", X"C8", X"E8", X"69", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"89", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"40", X"AD", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"89", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"40", X"40", X"8D", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"CD", X"C8", X"A8", X"00", X"00", X"00", X"C8", X"E8", X"64", X"A8", X"E8", X"40", X"00", X"00", X"20", X"E8", X"C8", X"49", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"AD", X"20", X"A4", X"00", X"00", X"00", X"64", X"40", X"84", X"64", X"40", X"84", X"00", X"00", X"20", X"64", X"60", X"D1", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"89", X"40", X"64", X"00", X"00", X"00", X"64", X"40", X"44", X"44", X"44", X"40", X"00", X"00", X"00", X"64", X"40", X"8D", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"AD", X"A8", X"84", X"00", X"00", X"00", X"A4", X"C8", X"44", X"A4", X"C8", X"20", X"00", X"00", X"20", X"C8", X"A4", X"49", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"CD", X"20", X"C8", X"00", X"00", X"00", X"84", X"44", X"C8", X"84", X"64", X"84", X"00", X"00", X"20", X"84", X"84", X"D1", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"92", X"44", X"60", X"20", X"48", X"69", X"69", X"64", X"40", X"44", X"69", X"69", X"49", X"44", X"20", X"64", X"69", X"B2", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"D1", X"C8", X"13", X"13", X"FB", X"A0", X"C4", X"D1", X"60", X"40", X"CD", X"C4", X"C8", X"CD", X"40", X"84", X"CC", X"C4", X"CC", X"A8", X"20", X"A8", X"C8", X"A4", X"C8", X"13", X"13", X"FA", X"A0", X"F6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"F1", X"CC", X"13", X"13", X"FB", X"C4", X"C8", X"D1", X"A4", X"A4", X"CD", X"C8", X"C8", X"CD", X"A4", X"A8", X"CC", X"C8", X"CC", X"A8", X"A4", X"A8", X"C8", X"C8", X"CC", X"13", X"13", X"FB", X"C4", X"FA", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"84", X"F1", X"B1", X"D1", X"40", X"20", X"AD", X"D1", X"CD", X"AD", X"40", X"40", X"CD", X"CD", X"F1", X"88", X"20", X"64", X"F1", X"AD", X"F1", X"64", X"20", X"88", X"F1", X"AD", X"D1", X"40", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"60", X"40", X"20", X"64", X"44", X"20", X"64", X"40", X"20", X"64", X"40", X"40", X"64", X"20", X"40", X"64", X"20", X"64", X"64", X"00", X"64", X"64", X"20", X"64", X"40", X"00", X"64", X"40", X"96", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"F5", X"64", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"E8", X"84", X"EC", X"C8", X"84", X"EC", X"A8", X"A8", X"EC", X"A4", X"C8", X"EC", X"84", X"C8", X"EC", X"84", X"C8", X"FA", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"60", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"44", X"40", X"00", X"00", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"40", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"60", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"40", X"00", X"00", X"00", X"00", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"40", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"F5", X"64", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"20", X"00", X"00", X"00", X"00", X"64", X"A8", X"A8", X"EC", X"A4", X"C8", X"EC", X"84", X"C8", X"EC", X"84", X"C8", X"FA", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"60", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"40", X"96", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"40", X"64", X"40", X"64", X"64", X"40", X"64", X"44", X"40", X"64", X"44", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"64", X"40", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"F5", X"60", X"C8", X"E8", X"40", X"C8", X"C8", X"40", X"C8", X"C8", X"64", X"C8", X"00", X"00", X"00", X"00", X"00", X"20", X"A4", X"84", X"E8", X"84", X"A4", X"E8", X"64", X"A8", X"E8", X"64", X"A4", X"FA", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"84", X"84", X"40", X"84", X"64", X"40", X"84", X"64", X"44", X"A4", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"60", X"96", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"40", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"44", X"44", X"44", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"40", X"64", X"64", X"40", X"44", X"64", X"40", X"44", X"40", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"D1", X"40", X"A4", X"C8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"00", X"00", X"00", X"00", X"00", X"20", X"84", X"84", X"C8", X"64", X"84", X"C8", X"64", X"84", X"C8", X"44", X"84", X"FA", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"D1", X"A4", X"84", X"44", X"C8", X"84", X"64", X"C8", X"84", X"64", X"C8", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"C8", X"84", X"B6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"B1", X"40", X"64", X"44", X"40", X"64", X"64", X"40", X"64", X"44", X"40", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"44", X"44", X"44", X"64", X"44", X"40", X"64", X"44", X"40", X"40", X"D6", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"D1", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"00", X"00", X"00", X"00", X"00", X"00", X"60", X"64", X"84", X"40", X"60", X"84", X"40", X"64", X"84", X"20", X"60", X"DB", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", X"13", 
X"CD", X"13", X"13", X"13", X"CD", X"CD", X"CD", X"13", X"13", X"13", X"CD", X"CD", X"F2", X"A8", X"64", X"F1", X"CD", X"CD", X"F1", X"A4", X"84", X"F1", X"CD", X"F1", X"F1", X"84", X"C8", X"F1", X"CD", X"D1", X"EC", X"40", X"EC", X"D1", X"CD", X"F1", X"C8", X"60", X"F1", X"CD", X"CD", X"F6", X"13", X"13", X"F6", X"CD", X"CD", X"13", X"13", X"13", X"CD", X"CD", X"CC", X"13", 
X"A4", X"13", X"13", X"13", X"C8", X"C8", X"C8", X"13", X"13", X"13", X"C4", X"C8", X"CD", X"40", X"40", X"AD", X"C8", X"C8", X"CD", X"40", X"40", X"CD", X"C4", X"C8", X"A9", X"40", X"64", X"CC", X"C8", X"CC", X"64", X"40", X"68", X"C8", X"C8", X"CC", X"64", X"40", X"A9", X"C8", X"C4", X"F1", X"13", X"13", X"F2", X"C4", X"A4", X"13", X"13", X"13", X"CC", X"C8", X"C4", X"13", 
X"40", X"13", X"13", X"13", X"88", X"60", X"44", X"13", X"13", X"13", X"64", X"60", X"8D", X"F1", X"F1", X"F6", X"40", X"40", X"D1", X"F1", X"F1", X"B1", X"40", X"44", X"D1", X"F1", X"F1", X"89", X"60", X"64", X"F1", X"F1", X"F2", X"64", X"60", X"89", X"F1", X"F1", X"D1", X"44", X"40", X"B2", X"13", X"13", X"B2", X"40", X"40", X"13", X"13", X"13", X"89", X"64", X"40", X"13", 
X"E8", X"C4", X"40", X"C4", X"E8", X"64", X"E8", X"C4", X"40", X"C4", X"E8", X"64", X"E8", X"A4", X"64", X"E8", X"C8", X"84", X"E8", X"A4", X"84", X"E8", X"A4", X"C8", X"E8", X"64", X"A4", X"E8", X"64", X"E8", X"E8", X"40", X"C8", X"E8", X"64", X"E8", X"C8", X"60", X"E8", X"C8", X"84", X"E8", X"80", X"84", X"E8", X"84", X"E8", X"C8", X"40", X"C4", X"E8", X"64", X"E8", X"C4", 
X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"40", X"64", X"40", X"40", X"64", X"20", X"44", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", 
X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"84", X"64", X"40", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"64", X"64", X"44", X"64", X"64", X"20", X"44", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", 
X"E8", X"EC", X"64", X"E8", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", X"EC", X"C8", X"A4", X"64", X"00", X"00", X"20", X"84", X"C8", X"EC", X"84", X"C8", X"EC", X"64", X"C8", X"00", X"00", X"00", X"84", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", X"EC", X"A4", X"A8", X"EC", X"64", X"E8", X"EC", X"64", X"E8", X"EC", X"64", X"EC", X"E8", 
X"64", X"20", X"64", X"64", X"20", X"64", X"40", X"20", X"64", X"20", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"64", X"20", X"64", X"44", X"20", X"84", X"00", X"00", X"00", X"00", X"00", X"64", X"20", X"44", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", 
X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"40", X"64", X"64", X"20", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"40", X"64", X"44", X"40", X"44", X"00", X"00", X"00", X"00", X"00", X"20", X"40", X"64", X"64", X"40", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", 
X"C8", X"E8", X"40", X"C8", X"C8", X"40", X"C8", X"C8", X"44", X"E8", X"C8", X"64", X"E8", X"A8", X"64", X"E8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"C8", X"E8", X"64", X"A8", X"E8", X"40", X"00", X"00", X"00", X"00", X"00", X"40", X"E8", X"C8", X"64", X"E8", X"A8", X"84", X"E8", X"84", X"A4", X"E8", X"64", X"C8", X"E8", X"64", X"C8", X"E8", X"44", X"C8", X"C8", 
X"84", X"20", X"84", X"84", X"20", X"A4", X"64", X"40", X"A4", X"44", X"64", X"A4", X"40", X"84", X"84", X"20", X"A4", X"20", X"00", X"00", X"00", X"00", X"00", X"64", X"40", X"84", X"64", X"40", X"84", X"00", X"00", X"00", X"00", X"00", X"20", X"44", X"64", X"84", X"40", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"A4", X"64", X"40", 
X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"44", X"44", X"44", X"44", X"44", X"40", X"64", X"44", X"40", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"40", X"44", X"44", X"44", X"40", X"00", X"00", X"00", X"00", X"00", X"20", X"44", X"64", X"44", X"40", X"64", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"40", 
X"A4", X"C8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"C8", X"84", X"44", X"C8", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"C8", X"44", X"A4", X"C8", X"20", X"00", X"00", X"00", X"00", X"00", X"40", X"C8", X"A8", X"40", X"C8", X"84", X"64", X"C8", X"64", X"84", X"C8", X"44", X"A4", X"C8", X"40", X"A8", X"C8", X"40", X"A8", X"A8", 
X"A8", X"40", X"C8", X"A8", X"40", X"C8", X"84", X"64", X"C8", X"64", X"84", X"C8", X"44", X"A4", X"C8", X"40", X"C8", X"20", X"00", X"00", X"00", X"00", X"00", X"84", X"44", X"C8", X"84", X"64", X"A4", X"00", X"00", X"00", X"00", X"00", X"40", X"64", X"84", X"C8", X"44", X"A4", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"C8", X"84", X"64", 
X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"44", X"40", X"64", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"20", X"64", X"64", X"40", X"44", X"44", X"44", X"44", X"44", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", 
X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"64", X"40", X"84", X"84", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"84", X"40", X"84", X"A4", X"20", X"00", X"00", X"00", X"00", X"00", X"20", X"84", X"84", X"20", X"84", X"64", X"40", X"A4", X"44", X"64", X"A4", X"40", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", 
X"C8", X"44", X"E8", X"C8", X"44", X"E8", X"A8", X"84", X"E8", X"84", X"A8", X"E8", X"64", X"C8", X"E8", X"40", X"E8", X"20", X"00", X"00", X"00", X"00", X"00", X"A8", X"64", X"E8", X"A8", X"84", X"C8", X"00", X"00", X"00", X"00", X"00", X"44", X"84", X"A8", X"E8", X"64", X"C8", X"E8", X"64", X"C8", X"C8", X"44", X"C8", X"C8", X"40", X"C8", X"C8", X"40", X"E8", X"A8", X"64", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"64", X"64", X"40", X"64", X"64", X"40", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"40", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"64", X"44", X"40", X"64", X"40", X"44", X"64", X"40", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"E8", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", X"EC", X"A4", X"C8", X"EC", X"84", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"E8", X"84", X"EC", X"C8", X"84", X"EC", X"A8", X"A8", X"EC", X"A4", X"C8", X"EC", X"84", X"C8", X"EC", X"84", X"E8", X"EC", X"64", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"20", X"64", X"40", X"40", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"E8", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", X"EC", X"A4", X"C8", X"EC", X"84", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"E8", X"84", X"EC", X"C8", X"A4", X"EC", X"A8", X"A8", X"EC", X"A4", X"C8", X"EC", X"84", X"C8", X"EC", X"84", X"E8", X"EC", X"64", X"E8", X"EC", X"64", X"EC", X"EC", X"64", X"EC", X"E8", X"64", X"EC", X"C8", X"84", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"00", X"00", X"20", X"64", X"20", X"64", X"40", X"40", X"64", X"40", X"44", X"40", X"00", X"00", X"40", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"00", X"00", X"00", X"64", X"20", X"64", X"40", X"40", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"00", X"00", X"00", X"00", X"20", X"44", X"64", X"44", X"40", X"64", X"40", X"40", X"00", X"00", X"00", X"00", X"20", X"64", X"64", X"20", X"64", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"44", X"64", X"40", X"44", X"64", X"40", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", 
X"C8", X"44", X"E8", X"C8", X"44", X"E8", X"A8", X"84", X"E8", X"84", X"A8", X"A8", X"00", X"00", X"00", X"00", X"00", X"C8", X"44", X"C8", X"C8", X"44", X"E8", X"20", X"00", X"00", X"00", X"00", X"44", X"A4", X"84", X"E8", X"84", X"A8", X"A8", X"00", X"00", X"00", X"00", X"00", X"C8", X"64", X"C8", X"C8", X"44", X"C8", X"C8", X"40", X"C8", X"C8", X"40", X"E8", X"A8", X"64", 
X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"84", X"64", X"44", X"A4", X"44", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"84", X"20", X"84", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"A4", X"44", X"64", X"A4", X"40", X"84", X"84", X"20", X"84", X"A4", X"20", X"84", X"84", 
X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"40", X"44", X"64", X"44", X"44", X"44", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"40", X"64", X"64", X"20", X"00", X"00", X"00", X"00", X"00", X"40", X"44", X"44", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", X"40", X"64", X"44", 
X"A8", X"40", X"C8", X"A8", X"40", X"C8", X"84", X"64", X"C8", X"64", X"84", X"64", X"00", X"00", X"00", X"00", X"00", X"84", X"40", X"A8", X"A8", X"40", X"A8", X"00", X"00", X"00", X"00", X"00", X"20", X"84", X"84", X"C8", X"64", X"84", X"64", X"00", X"00", X"00", X"00", X"00", X"84", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"C8", X"84", X"64", 
X"A4", X"C8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"40", X"A8", X"A8", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"C8", X"84", X"64", X"C8", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"A8", X"A8", X"40", X"A8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"C8", X"64", X"84", X"C8", X"44", X"A4", X"C8", X"40", X"A8", X"C8", X"40", X"A8", X"A8", 
X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"44", X"44", X"44", X"64", X"20", X"00", X"00", X"00", X"00", X"00", X"40", X"40", X"64", X"44", X"40", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"44", X"44", X"44", X"64", X"20", X"00", X"00", X"00", X"00", X"00", X"40", X"40", X"44", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"40", X"44", X"64", X"40", 
X"84", X"20", X"84", X"84", X"20", X"A4", X"64", X"40", X"A4", X"44", X"64", X"44", X"00", X"00", X"00", X"00", X"00", X"64", X"20", X"84", X"84", X"20", X"84", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"84", X"44", X"64", X"64", X"00", X"00", X"00", X"00", X"00", X"64", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"A4", X"64", X"40", 
X"C8", X"E8", X"40", X"C8", X"C8", X"40", X"C8", X"C8", X"44", X"E8", X"C8", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"E8", X"A4", X"84", X"E8", X"84", X"00", X"00", X"00", X"00", X"00", X"20", X"C8", X"C8", X"40", X"C8", X"E8", X"00", X"00", X"00", X"00", X"00", X"00", X"84", X"E8", X"84", X"A4", X"E8", X"64", X"C8", X"E8", X"64", X"C8", X"E8", X"44", X"C8", X"C8", 
X"64", X"20", X"64", X"64", X"20", X"64", X"44", X"40", X"64", X"40", X"64", X"20", X"00", X"00", X"00", X"00", X"00", X"44", X"20", X"64", X"64", X"20", X"64", X"00", X"00", X"00", X"00", X"00", X"00", X"44", X"44", X"64", X"40", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"40", X"40", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"20", X"64", X"64", X"40", 
X"84", X"20", X"84", X"84", X"40", X"84", X"64", X"44", X"84", X"44", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"64", X"20", X"84", X"64", X"40", X"84", X"00", X"00", X"00", X"00", X"00", X"00", X"64", X"64", X"84", X"44", X"64", X"40", X"00", X"00", X"00", X"00", X"00", X"64", X"40", X"64", X"84", X"20", X"84", X"84", X"20", X"84", X"84", X"20", X"84", X"64", X"40"



);
begin

	Q <= castle(ADDR);		
			
end arch;
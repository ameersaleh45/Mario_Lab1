--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity coin_sound is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(12 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end coin_sound;

architecture arch of coin_sound is

type table_type is array(0 to 8191) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FD",
X"FB",
X"FC",
X"00",
X"02",
X"04",
X"07",
X"05",
X"04",
X"02",
X"FD",
X"FA",
X"FA",
X"FA",
X"FE",
X"01",
X"05",
X"09",
X"08",
X"05",
X"02",
X"FD",
X"F7",
X"F7",
X"F7",
X"FD",
X"02",
X"06",
X"0B",
X"0A",
X"06",
X"03",
X"FD",
X"F6",
X"F5",
X"F5",
X"FA",
X"02",
X"08",
X"0C",
X"0D",
X"08",
X"02",
X"FD",
X"F4",
X"F2",
X"F4",
X"F9",
X"01",
X"08",
X"0D",
X"0E",
X"09",
X"04",
X"FF",
X"F4",
X"F1",
X"F3",
X"F7",
X"00",
X"09",
X"0C",
X"10",
X"0C",
X"03",
X"FE",
X"F5",
X"EF",
X"F1",
X"F5",
X"FE",
X"08",
X"0D",
X"0F",
X"0D",
X"06",
X"FF",
X"F4",
X"EF",
X"EF",
X"F4",
X"FC",
X"05",
X"0D",
X"10",
X"0F",
X"08",
X"FF",
X"F6",
X"EE",
X"ED",
X"F3",
X"FA",
X"05",
X"0E",
X"10",
X"11",
X"0B",
X"01",
X"F8",
X"EF",
X"EC",
X"F0",
X"F7",
X"02",
X"0D",
X"11",
X"12",
X"0D",
X"02",
X"FA",
X"F1",
X"ED",
X"F0",
X"F6",
X"00",
X"0A",
X"0F",
X"11",
X"0D",
X"04",
X"FC",
X"F4",
X"F0",
X"F1",
X"F6",
X"FF",
X"07",
X"0D",
X"0E",
X"0C",
X"05",
X"FE",
X"F7",
X"F2",
X"F2",
X"F6",
X"FD",
X"04",
X"0B",
X"0D",
X"0B",
X"06",
X"FF",
X"F9",
X"F4",
X"F3",
X"F7",
X"FD",
X"03",
X"09",
X"0B",
X"0A",
X"06",
X"00",
X"FA",
X"F6",
X"F5",
X"F7",
X"FD",
X"02",
X"07",
X"0A",
X"0A",
X"06",
X"00",
X"FB",
X"F7",
X"F6",
X"F7",
X"FC",
X"01",
X"06",
X"09",
X"09",
X"06",
X"01",
X"FC",
X"F8",
X"F7",
X"F8",
X"FC",
X"01",
X"05",
X"09",
X"09",
X"06",
X"01",
X"FC",
X"F8",
X"F7",
X"F8",
X"FC",
X"01",
X"05",
X"08",
X"08",
X"06",
X"01",
X"FD",
X"F9",
X"F7",
X"F9",
X"FC",
X"00",
X"05",
X"08",
X"08",
X"06",
X"01",
X"FD",
X"F9",
X"F8",
X"F9",
X"FC",
X"00",
X"04",
X"07",
X"08",
X"06",
X"02",
X"FE",
X"FA",
X"F8",
X"F9",
X"FB",
X"00",
X"04",
X"07",
X"08",
X"06",
X"02",
X"FF",
X"FB",
X"F8",
X"F9",
X"FB",
X"00",
X"03",
X"06",
X"07",
X"06",
X"03",
X"FF",
X"FC",
X"F9",
X"FA",
X"FC",
X"00",
X"03",
X"07",
X"08",
X"07",
X"04",
X"00",
X"FC",
X"FA",
X"F9",
X"FB",
X"FF",
X"02",
X"05",
X"07",
X"06",
X"04",
X"00",
X"FD",
X"FA",
X"FA",
X"FB",
X"FF",
X"02",
X"05",
X"07",
X"07",
X"04",
X"01",
X"FE",
X"FB",
X"F9",
X"FB",
X"FE",
X"01",
X"04",
X"06",
X"06",
X"04",
X"01",
X"FE",
X"FB",
X"FA",
X"FB",
X"FE",
X"01",
X"04",
X"06",
X"07",
X"05",
X"02",
X"FF",
X"FC",
X"FA",
X"FA",
X"FD",
X"00",
X"03",
X"05",
X"06",
X"05",
X"01",
X"FF",
X"FC",
X"FA",
X"FB",
X"FD",
X"00",
X"03",
X"06",
X"06",
X"05",
X"02",
X"00",
X"FD",
X"FB",
X"FB",
X"FC",
X"00",
X"02",
X"04",
X"05",
X"05",
X"02",
X"00",
X"FD",
X"FB",
X"FB",
X"FD",
X"00",
X"02",
X"05",
X"06",
X"05",
X"03",
X"00",
X"FE",
X"FB",
X"FB",
X"FC",
X"FF",
X"01",
X"04",
X"05",
X"05",
X"03",
X"00",
X"FE",
X"FC",
X"FB",
X"FD",
X"FF",
X"01",
X"04",
X"05",
X"05",
X"03",
X"01",
X"FF",
X"FC",
X"FB",
X"FC",
X"FE",
X"00",
X"03",
X"04",
X"04",
X"03",
X"01",
X"FF",
X"FC",
X"FC",
X"FC",
X"FE",
X"00",
X"03",
X"05",
X"05",
X"04",
X"01",
X"FF",
X"FD",
X"FC",
X"FC",
X"FE",
X"00",
X"02",
X"04",
X"04",
X"03",
X"01",
X"FF",
X"FD",
X"FC",
X"FC",
X"FE",
X"00",
X"02",
X"04",
X"05",
X"04",
X"02",
X"00",
X"FE",
X"FC",
X"FC",
X"FD",
X"00",
X"01",
X"03",
X"04",
X"03",
X"02",
X"00",
X"FE",
X"FC",
X"FC",
X"FE",
X"00",
X"01",
X"03",
X"04",
X"04",
X"02",
X"00",
X"FF",
X"FD",
X"FC",
X"FD",
X"FF",
X"00",
X"02",
X"03",
X"03",
X"02",
X"00",
X"FF",
X"FD",
X"FD",
X"FD",
X"FF",
X"01",
X"03",
X"04",
X"04",
X"03",
X"00",
X"FF",
X"FD",
X"FD",
X"FD",
X"FF",
X"00",
X"02",
X"03",
X"03",
X"02",
X"00",
X"FF",
X"FE",
X"FD",
X"FD",
X"FF",
X"00",
X"02",
X"03",
X"04",
X"03",
X"01",
X"00",
X"FE",
X"FD",
X"FD",
X"FE",
X"00",
X"01",
X"03",
X"03",
X"03",
X"01",
X"00",
X"FE",
X"FD",
X"FD",
X"FE",
X"00",
X"01",
X"03",
X"03",
X"03",
X"01",
X"00",
X"FF",
X"FD",
X"FD",
X"FE",
X"00",
X"01",
X"02",
X"03",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FD",
X"FE",
X"00",
X"01",
X"02",
X"03",
X"03",
X"02",
X"00",
X"FF",
X"FE",
X"FD",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"02",
X"00",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"00",
X"02",
X"03",
X"03",
X"02",
X"00",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"02",
X"00",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"03",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FE",
X"FE",
X"FF",
X"00",
X"01",
X"01",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"01",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FD",
X"FE",
X"01",
X"04",
X"04",
X"03",
X"02",
X"FC",
X"FB",
X"FD",
X"FF",
X"04",
X"07",
X"05",
X"02",
X"FE",
X"F9",
X"F9",
X"FE",
X"03",
X"07",
X"07",
X"05",
X"FE",
X"F8",
X"F8",
X"FA",
X"01",
X"09",
X"09",
X"05",
X"01",
X"F8",
X"F4",
X"F9",
X"FF",
X"07",
X"0B",
X"08",
X"02",
X"FB",
X"F5",
X"F6",
X"FD",
X"06",
X"0B",
X"0A",
X"04",
X"FD",
X"F4",
X"F4",
X"FA",
X"01",
X"0A",
X"0B",
X"06",
X"00",
X"F6",
X"F2",
X"F7",
X"00",
X"07",
X"0C",
X"0A",
X"02",
X"F8",
X"F2",
X"F4",
X"FB",
X"06",
X"0D",
X"0C",
X"07",
X"FE",
X"F3",
X"F1",
X"F7",
X"01",
X"0B",
X"0E",
X"09",
X"00",
X"F7",
X"F1",
X"F4",
X"FE",
X"07",
X"0D",
X"0C",
X"04",
X"FA",
X"F3",
X"F3",
X"FA",
X"04",
X"0C",
X"0D",
X"07",
X"FE",
X"F5",
X"F2",
X"F7",
X"00",
X"09",
X"0E",
X"0A",
X"00",
X"F7",
X"F2",
X"F4",
X"FD",
X"06",
X"0D",
X"0B",
X"04",
X"FB",
X"F4",
X"F4",
X"FB",
X"03",
X"0B",
X"0C",
X"06",
X"FE",
X"F7",
X"F4",
X"F8",
X"00",
X"08",
X"0B",
X"08",
X"00",
X"F9",
X"F5",
X"F7",
X"FF",
X"06",
X"0A",
X"09",
X"02",
X"FA",
X"F5",
X"F6",
X"FC",
X"04",
X"09",
X"09",
X"04",
X"FD",
X"F7",
X"F6",
X"FB",
X"02",
X"08",
X"0A",
X"06",
X"FF",
X"F8",
X"F6",
X"F9",
X"00",
X"06",
X"09",
X"07",
X"01",
X"FB",
X"F6",
X"F8",
X"FE",
X"04",
X"09",
X"09",
X"03",
X"FD",
X"F7",
X"F7",
X"FC",
X"02",
X"08",
X"09",
X"05",
X"FF",
X"F9",
X"F7",
X"FB",
X"01",
X"07",
X"0A",
X"08",
X"01",
X"FB",
X"F7",
X"F8",
X"FF",
X"04",
X"08",
X"08",
X"03",
X"FD",
X"F8",
X"F9",
X"FD",
X"03",
X"08",
X"09",
X"05",
X"00",
X"FA",
X"F7",
X"FB",
X"00",
X"05",
X"08",
X"06",
X"00",
X"FB",
X"F8",
X"FA",
X"FF",
X"05",
X"09",
X"08",
X"03",
X"FE",
X"F9",
X"F8",
X"FD",
X"02",
X"06",
X"08",
X"04",
X"FF",
X"FA",
X"F9",
X"FC",
X"01",
X"06",
X"08",
X"06",
X"01",
X"FC",
X"F9",
X"FA",
X"FF",
X"04",
X"07",
X"06",
X"02",
X"FD",
X"FA",
X"FA",
X"FE",
X"03",
X"07",
X"08",
X"05",
X"00",
X"FB",
X"F9",
X"FB",
X"00",
X"05",
X"07",
X"05",
X"00",
X"FC",
X"F9",
X"FB",
X"00",
X"04",
X"07",
X"07",
X"02",
X"FE",
X"FA",
X"F9",
X"FD",
X"02",
X"05",
X"06",
X"03",
X"FF",
X"FB",
X"FA",
X"FC",
X"00",
X"05",
X"07",
X"05",
X"01",
X"FD",
X"FA",
X"FB",
X"FF",
X"03",
X"06",
X"06",
X"02",
X"FE",
X"FB",
X"FB",
X"FE",
X"02",
X"06",
X"06",
X"04",
X"00",
X"FC",
X"FA",
X"FC",
X"00",
X"04",
X"06",
X"04",
X"00",
X"FD",
X"FA",
X"FC",
X"00",
X"04",
X"06",
X"06",
X"02",
X"FE",
X"FB",
X"FB",
X"FE",
X"01",
X"05",
X"05",
X"03",
X"FF",
X"FC",
X"FB",
X"FD",
X"01",
X"04",
X"06",
X"04",
X"00",
X"FD",
X"FB",
X"FC",
X"FF",
X"03",
X"05",
X"05",
X"01",
X"FE",
X"FB",
X"FC",
X"FF",
X"02",
X"05",
X"06",
X"03",
X"00",
X"FC",
X"FB",
X"FD",
X"00",
X"03",
X"05",
X"04",
X"00",
X"FD",
X"FB",
X"FD",
X"00",
X"03",
X"05",
X"05",
X"02",
X"FF",
X"FC",
X"FC",
X"FE",
X"01",
X"04",
X"04",
X"02",
X"FF",
X"FC",
X"FC",
X"FE",
X"00",
X"04",
X"05",
X"04",
X"00",
X"FE",
X"FC",
X"FC",
X"00",
X"02",
X"04",
X"04",
X"01",
X"FE",
X"FC",
X"FC",
X"FF",
X"02",
X"04",
X"05",
X"02",
X"00",
X"FD",
X"FC",
X"FD",
X"00",
X"03",
X"04",
X"03",
X"00",
X"FE",
X"FC",
X"FD",
X"00",
X"02",
X"04",
X"04",
X"01",
X"FF",
X"FC",
X"FC",
X"FF",
X"01",
X"03",
X"04",
X"02",
X"00",
X"FD",
X"FC",
X"FE",
X"00",
X"03",
X"04",
X"03",
X"00",
X"FE",
X"FC",
X"FD",
X"00",
X"02",
X"03",
X"03",
X"01",
X"FF",
X"FD",
X"FD",
X"FF",
X"01",
X"04",
X"04",
X"02",
X"00",
X"FD",
X"FC",
X"FE",
X"00",
X"02",
X"03",
X"02",
X"00",
X"FE",
X"FD",
X"FE",
X"00",
X"02",
X"04",
X"03",
X"01",
X"FF",
X"FD",
X"FD",
X"FF",
X"01",
X"03",
X"03",
X"01",
X"00",
X"FD",
X"FD",
X"FF",
X"00",
X"03",
X"04",
X"02",
X"00",
X"FE",
X"FD",
X"FE",
X"00",
X"01",
X"03",
X"03",
X"00",
X"FF",
X"FD",
X"FE",
X"00",
X"01",
X"03",
X"03",
X"01",
X"00",
X"FE",
X"FD",
X"FE",
X"00",
X"02",
X"03",
X"02",
X"00",
X"FE",
X"FD",
X"FE",
X"00",
X"02",
X"03",
X"03",
X"01",
X"FF",
X"FE",
X"FE",
X"FF",
X"01",
X"02",
X"02",
X"01",
X"00",
X"FE",
X"FE",
X"FF",
X"00",
X"02",
X"03",
X"02",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"01",
X"02",
X"02",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"01",
X"02",
X"03",
X"01",
X"00",
X"FE",
X"FE",
X"FF",
X"00",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"00",
X"02",
X"02",
X"01",
X"00",
X"FE",
X"FE",
X"FF",
X"00",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"01",
X"02",
X"02",
X"00",
X"FF",
X"FE",
X"FE",
X"00",
X"01",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"02",
X"00",
X"00",
X"FE",
X"FE",
X"00",
X"00",
X"01",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"01",
X"02",
X"01",
X"00",
X"FF",
X"FE",
X"FF",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"02",
X"02",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"02",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"


);

begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;
--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Small_mario_jump_sound is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(13 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end Small_mario_jump_sound;

architecture arch of Small_mario_jump_sound is

type table_type is array(0 to 16383) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"06",
X"1F",
X"1D",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"11",
X"F7",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"14",
X"18",
X"17",
X"16",
X"16",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"13",
X"14",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"0F",
X"11",
X"F8",
X"F0",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F4",
X"F8",
X"F3",
X"0F",
X"1F",
X"1A",
X"1C",
X"1A",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"16",
X"16",
X"15",
X"16",
X"14",
X"15",
X"13",
X"15",
X"12",
X"16",
X"00",
X"E9",
X"EF",
X"EC",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F1",
X"F3",
X"F1",
X"F4",
X"F0",
X"00",
X"1C",
X"17",
X"19",
X"17",
X"18",
X"16",
X"17",
X"16",
X"16",
X"15",
X"16",
X"14",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"10",
X"13",
X"06",
X"E8",
X"EC",
X"EA",
X"EC",
X"EB",
X"ED",
X"EC",
X"ED",
X"EC",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F5",
X"16",
X"17",
X"17",
X"16",
X"17",
X"15",
X"16",
X"15",
X"15",
X"14",
X"15",
X"13",
X"14",
X"13",
X"13",
X"12",
X"13",
X"11",
X"12",
X"11",
X"12",
X"10",
X"11",
X"0F",
X"11",
X"F2",
X"E8",
X"EB",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EE",
X"F0",
X"EF",
X"F1",
X"EF",
X"F2",
X"ED",
X"06",
X"1A",
X"15",
X"17",
X"15",
X"16",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"11",
X"0E",
X"12",
X"01",
X"E6",
X"EB",
X"E8",
X"EB",
X"EA",
X"EB",
X"EB",
X"EC",
X"EB",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"EF",
X"F6",
X"17",
X"16",
X"17",
X"15",
X"16",
X"14",
X"15",
X"14",
X"14",
X"13",
X"14",
X"12",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"EF",
X"E8",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EE",
X"F0",
X"EE",
X"F2",
X"ED",
X"08",
X"19",
X"15",
X"17",
X"15",
X"15",
X"14",
X"13",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0D",
X"0F",
X"0C",
X"10",
X"00",
X"E6",
X"EB",
X"E9",
X"EB",
X"EA",
X"EC",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F1",
X"EF",
X"F8",
X"15",
X"13",
X"14",
X"13",
X"14",
X"12",
X"13",
X"11",
X"12",
X"11",
X"12",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0C",
X"EE",
X"E9",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"F0",
X"EF",
X"F0",
X"EF",
X"F1",
X"EF",
X"F2",
X"EE",
X"09",
X"17",
X"13",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0E",
X"0F",
X"0E",
X"0F",
X"0C",
X"11",
X"FE",
X"E7",
X"EC",
X"EA",
X"EC",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F2",
X"EF",
X"FA",
X"16",
X"13",
X"15",
X"13",
X"14",
X"12",
X"13",
X"12",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0B",
X"ED",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"EF",
X"F1",
X"F0",
X"F2",
X"EF",
X"0C",
X"17",
X"13",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"10",
X"0E",
X"10",
X"0C",
X"11",
X"FC",
X"E7",
X"EC",
X"EA",
X"EC",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F2",
X"EF",
X"FC",
X"17",
X"13",
X"15",
X"13",
X"14",
X"12",
X"13",
X"12",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0F",
X"0A",
X"EB",
X"EB",
X"EA",
X"EC",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F2",
X"F0",
X"0C",
X"13",
X"11",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0E",
X"0C",
X"0E",
X"0B",
X"0F",
X"F9",
X"E8",
X"ED",
X"EB",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F1",
X"F0",
X"F2",
X"F0",
X"F3",
X"EF",
X"FE",
X"15",
X"11",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0C",
X"0E",
X"07",
X"EB",
X"EC",
X"EB",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F1",
X"F0",
X"F2",
X"F1",
X"F3",
X"F1",
X"0B",
X"14",
X"12",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0D",
X"0E",
X"0D",
X"0E",
X"0B",
X"10",
X"FE",
X"E9",
X"EE",
X"EB",
X"ED",
X"EC",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F1",
X"F7",
X"13",
X"12",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0E",
X"0F",
X"0E",
X"0F",
X"0D",
X"0E",
X"0D",
X"0E",
X"0C",
X"0E",
X"F4",
X"EA",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F1",
X"F1",
X"F2",
X"F1",
X"F3",
X"EF",
X"00",
X"16",
X"11",
X"14",
X"11",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0E",
X"07",
X"EC",
X"ED",
X"EC",
X"ED",
X"EC",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F2",
X"F1",
X"F2",
X"F1",
X"F3",
X"F1",
X"0B",
X"15",
X"0F",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0D",
X"0B",
X"0C",
X"0B",
X"0C",
X"0A",
X"0E",
X"FE",
X"EA",
X"EE",
X"EC",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F3",
X"F2",
X"F8",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0C",
X"0B",
X"0C",
X"F4",
X"EC",
X"EE",
X"ED",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F1",
X"F2",
X"F2",
X"F3",
X"F2",
X"F4",
X"F0",
X"00",
X"14",
X"10",
X"12",
X"10",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0B",
X"0D",
X"07",
X"ED",
X"EE",
X"ED",
X"EF",
X"EE",
X"EF",
X"EE",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F1",
X"F1",
X"F2",
X"F1",
X"F2",
X"F1",
X"F3",
X"F2",
X"F3",
X"F2",
X"F4",
X"F2",
X"0B",
X"13",
X"10",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"0A",
X"0E",
X"FF",
X"EB",
X"EF",
X"ED",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F2",
X"F4",
X"F2",
X"FA",
X"19",
X"19",
X"19",
X"18",
X"18",
X"18",
X"17",
X"17",
X"16",
X"17",
X"14",
X"18",
X"03",
X"EB",
X"F1",
X"EE",
X"F1",
X"EF",
X"F1",
X"F0",
X"F1",
X"F0",
X"F2",
X"F1",
X"F2",
X"F1",
X"F3",
X"F2",
X"F3",
X"F2",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F5",
X"F8",
X"F3",
X"07",
X"20",
X"1B",
X"1D",
X"1B",
X"1B",
X"1A",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"19",
X"FB",
X"EF",
X"F3",
X"F1",
X"F3",
X"F2",
X"F3",
X"F2",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"15",
X"20",
X"1C",
X"1E",
X"1C",
X"1C",
X"1B",
X"1C",
X"1A",
X"1B",
X"19",
X"1B",
X"12",
X"F2",
X"F3",
X"F2",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F7",
X"FF",
X"1E",
X"1E",
X"1E",
X"1D",
X"1D",
X"1D",
X"1B",
X"1C",
X"1A",
X"1C",
X"18",
X"1D",
X"07",
X"F0",
X"F5",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FB",
X"1B",
X"20",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"1A",
X"1C",
X"13",
X"F4",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"0C",
X"22",
X"1D",
X"1F",
X"1D",
X"1D",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"19",
X"1C",
X"00",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FE",
X"1D",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"19",
X"1C",
X"11",
X"F2",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"10",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1B",
X"FF",
X"F1",
X"F5",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FA",
X"F7",
X"00",
X"1F",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"0E",
X"F1",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"13",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1B",
X"1B",
X"1B",
X"1A",
X"1A",
X"FB",
X"F1",
X"F5",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"02",
X"21",
X"1E",
X"1F",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"0A",
X"F0",
X"F5",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"16",
X"21",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1B",
X"18",
X"F9",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"05",
X"21",
X"1E",
X"1F",
X"1D",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"07",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"19",
X"21",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1B",
X"16",
X"F6",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"09",
X"22",
X"1D",
X"1F",
X"1D",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"03",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FC",
X"1B",
X"20",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1C",
X"14",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"0C",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1C",
X"00",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FE",
X"1D",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"19",
X"1C",
X"11",
X"F2",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"10",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1B",
X"FE",
X"F1",
X"F5",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FA",
X"F7",
X"00",
X"1F",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"0E",
X"F1",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"13",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1B",
X"1B",
X"1B",
X"1A",
X"1A",
X"FB",
X"F1",
X"F5",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"02",
X"21",
X"1E",
X"1F",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"0A",
X"F0",
X"F5",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"16",
X"21",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1B",
X"18",
X"F9",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"05",
X"21",
X"1E",
X"1F",
X"1D",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"07",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"19",
X"21",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1B",
X"16",
X"F6",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"09",
X"22",
X"1D",
X"1F",
X"1D",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"03",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FC",
X"1B",
X"20",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"1A",
X"1C",
X"14",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"FB",
X"F6",
X"0C",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1C",
X"00",
X"F0",
X"F6",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FE",
X"1D",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"19",
X"1C",
X"11",
X"F2",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"10",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1B",
X"FE",
X"F1",
X"F5",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FA",
X"F7",
X"00",
X"1F",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1D",
X"1B",
X"1C",
X"19",
X"1D",
X"0D",
X"F1",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F7",
X"13",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1A",
X"FB",
X"F1",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"00",
X"1F",
X"1E",
X"1F",
X"1E",
X"1E",
X"1D",
X"1C",
X"1C",
X"1B",
X"1B",
X"1A",
X"1B",
X"15",
X"F4",
X"F4",
X"F3",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"FA",
X"1A",
X"20",
X"1E",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1B",
X"19",
X"1A",
X"FB",
X"F2",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"12",
X"22",
X"1D",
X"1F",
X"1D",
X"1D",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"02",
X"F0",
X"F5",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F8",
X"FB",
X"F6",
X"08",
X"22",
X"1D",
X"1F",
X"1D",
X"1E",
X"1D",
X"1C",
X"1C",
X"1B",
X"1C",
X"19",
X"1D",
X"0B",
X"F0",
X"F5",
X"F2",
X"F5",
X"F3",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F8",
X"FE",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0B",
X"F6",
X"F6",
X"F5",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"11",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"FB",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FC",
X"FA",
X"FC",
X"F9",
X"0C",
X"15",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"12",
X"10",
X"12",
X"00",
X"F5",
X"F9",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FC",
X"FA",
X"FD",
X"F9",
X"05",
X"16",
X"13",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"12",
X"10",
X"13",
X"06",
X"F5",
X"F9",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FA",
X"00",
X"15",
X"13",
X"14",
X"13",
X"13",
X"12",
X"13",
X"12",
X"12",
X"12",
X"11",
X"12",
X"0C",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FD",
X"12",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"11",
X"FB",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"0D",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"13",
X"00",
X"F6",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"FD",
X"F9",
X"07",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"13",
X"06",
X"F5",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"00",
X"16",
X"13",
X"14",
X"13",
X"13",
X"12",
X"13",
X"12",
X"12",
X"12",
X"11",
X"12",
X"0C",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FD",
X"13",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"10",
X"FB",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"0E",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"12",
X"00",
X"F6",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"FD",
X"F9",
X"07",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"13",
X"05",
X"F5",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"01",
X"16",
X"13",
X"14",
X"13",
X"13",
X"12",
X"13",
X"12",
X"12",
X"12",
X"11",
X"12",
X"0B",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FB",
X"FE",
X"13",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"11",
X"10",
X"FA",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"0E",
X"15",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"12",
X"00",
X"F6",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"FD",
X"F9",
X"08",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"12",
X"10",
X"13",
X"04",
X"F5",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"02",
X"16",
X"13",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"12",
X"0A",
X"F6",
X"F9",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FE",
X"13",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"FE",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"00",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"10",
X"FB",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"01",
X"16",
X"13",
X"14",
X"13",
X"13",
X"12",
X"13",
X"12",
X"12",
X"11",
X"12",
X"0E",
X"F9",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"03",
X"16",
X"13",
X"14",
X"13",
X"14",
X"12",
X"13",
X"11",
X"12",
X"11",
X"12",
X"0C",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"F9",
X"06",
X"17",
X"12",
X"15",
X"12",
X"14",
X"12",
X"13",
X"11",
X"13",
X"10",
X"13",
X"09",
X"F7",
X"F9",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"09",
X"17",
X"12",
X"15",
X"12",
X"14",
X"12",
X"13",
X"11",
X"13",
X"10",
X"13",
X"07",
X"F6",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FA",
X"0A",
X"13",
X"10",
X"12",
X"10",
X"11",
X"0F",
X"11",
X"0F",
X"10",
X"0E",
X"11",
X"03",
X"F6",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"0C",
X"13",
X"10",
X"12",
X"10",
X"11",
X"10",
X"11",
X"0F",
X"10",
X"0E",
X"11",
X"01",
X"F7",
X"FA",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"0F",
X"13",
X"11",
X"12",
X"10",
X"11",
X"10",
X"11",
X"0F",
X"10",
X"0E",
X"11",
X"00",
X"F7",
X"FA",
X"F8",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FB",
X"FE",
X"11",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0F",
X"10",
X"FE",
X"F7",
X"FA",
X"F8",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"00",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0E",
X"FC",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"00",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0D",
X"FA",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"02",
X"14",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0B",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"05",
X"14",
X"11",
X"12",
X"10",
X"11",
X"10",
X"11",
X"0F",
X"10",
X"0E",
X"11",
X"09",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"07",
X"14",
X"10",
X"12",
X"10",
X"12",
X"10",
X"11",
X"0F",
X"11",
X"0E",
X"11",
X"06",
X"F7",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"0A",
X"14",
X"11",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"11",
X"09",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"0F",
X"12",
X"11",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"11",
X"03",
X"F7",
X"FA",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"00",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"FF",
X"F7",
X"FA",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"05",
X"14",
X"11",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"10",
X"0D",
X"FA",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"0B",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"11",
X"08",
X"F7",
X"FA",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"10",
X"12",
X"11",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"11",
X"02",
X"F7",
X"FA",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"00",
X"13",
X"11",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"FE",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"06",
X"14",
X"11",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"10",
X"0C",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"0A",
X"10",
X"0E",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0E",
X"06",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FE",
X"0F",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0F",
X"00",
X"F8",
X"FB",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"FB",
X"FD",
X"FB",
X"01",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"FD",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"FD",
X"FA",
X"07",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"0A",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"0C",
X"11",
X"0F",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0D",
X"0F",
X"05",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"0F",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0F",
X"00",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"02",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"FC",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"08",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"09",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"0C",
X"11",
X"0F",
X"10",
X"0E",
X"0F",
X"0E",
X"0F",
X"0D",
X"0F",
X"09",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"0F",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0D",
X"0F",
X"05",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"FB",
X"FD",
X"FB",
X"01",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0D",
X"0F",
X"00",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"FD",
X"FA",
X"06",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"FE",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"0A",
X"11",
X"0F",
X"10",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0E",
X"0B",
X"FB",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FE",
X"0E",
X"10",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0F",
X"0D",
X"0F",
X"07",
X"F9",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0D",
X"0F",
X"03",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"FD",
X"FA",
X"03",
X"11",
X"0F",
X"10",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0D",
X"0E",
X"00",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"FD",
X"FB",
X"08",
X"11",
X"0F",
X"10",
X"0E",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"FC",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"0C",
X"11",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0F",
X"09",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"0F",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0F",
X"0D",
X"0F",
X"05",
X"F8",
X"FB",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"0E",
X"0C",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"00",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FB",
X"04",
X"0F",
X"0C",
X"0D",
X"0C",
X"0D",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"FE",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"08",
X"0F",
X"0C",
X"0D",
X"0C",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"09",
X"FC",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"0C",
X"0E",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0C",
X"0B",
X"0D",
X"06",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0B",
X"0D",
X"03",
X"F9",
X"FC",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"FB",
X"02",
X"0F",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0B",
X"0D",
X"00",
X"F9",
X"FC",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"FB",
X"06",
X"0F",
X"0C",
X"0E",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"06",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0E",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"07",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0E",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"07",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0E",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"07",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"08",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0D",
X"0B",
X"0D",
X"08",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0D",
X"08",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0C",
X"09",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"09",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"09",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FF",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"09",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FF",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0A",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FE",
X"0C",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0A",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FC",
X"FE",
X"0C",
X"0E",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0A",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"08",
X"FC",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"0A",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"09",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"09",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"09",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"09",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"FE",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"FF",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"07",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0B",
X"04",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"08",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0B",
X"03",
X"FA",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"01",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"09",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"09",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"09",
X"0B",
X"02",
X"FA",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"02",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"08",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"0A",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"09",
X"0B",
X"00",
X"FA",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"04",
X"0C",
X"0A",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"07",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FF",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0B",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"05",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0B",
X"06",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"00",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"06",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0B",
X"05",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"FE",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"07",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0B",
X"03",
X"FA",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"00",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"09",
X"FD",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"09",
X"0C",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"09",
X"0B",
X"02",
X"FA",
X"FD",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FC",
X"01",
X"0A",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"06",
X"FD",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"07",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"09",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"02",
X"0A",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"09",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FC",
X"01",
X"0A",
X"08",
X"09",
X"09",
X"08",
X"08",
X"08",
X"09",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"0A",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"01",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"02",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"03",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"08",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"04",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"07",
X"0A",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"05",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"07",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"09",
X"06",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"06",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"07",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"05",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"08",
X"FF",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"03",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"08",
X"00",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"02",
X"0A",
X"08",
X"09",
X"09",
X"08",
X"08",
X"08",
X"09",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"01",
X"0A",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"0A",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"01",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"02",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"00",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"03",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FF",
X"08",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"04",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"07",
X"0A",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"06",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"06",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"09",
X"06",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"05",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"07",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"04",
X"0A",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"08",
X"FF",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"02",
X"07",
X"06",
X"07",
X"06",
X"06",
X"05",
X"07",
X"01",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"04",
X"07",
X"06",
X"07",
X"06",
X"07",
X"05",
X"07",
X"00",
X"FC",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"06",
X"FF",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FD",
X"00",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"04",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"03",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"01",
X"FC",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"05",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FD",
X"01",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"03",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"04",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"06",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"06",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"04",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"02",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"02",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"05",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"07",
X"07",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FD",
X"00",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"04",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"03",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"01",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"06",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"07",
X"05",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FD",
X"01",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"03",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"04",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"06",
X"07",
X"07",
X"07",
X"06",
X"06",
X"06",
X"06",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"00",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"04",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"02",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"02",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"07",
X"06",
X"07",
X"06",
X"07",
X"06",
X"07",
X"00",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"03",
X"08",
X"06",
X"07",
X"06",
X"07",
X"06",
X"05",
X"FE",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"07",
X"01",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"01",
X"05",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"05",
X"01",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"04",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"04",
X"05",
X"05",
X"04",
X"04",
X"04",
X"05",
X"02",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"03",
X"05",
X"04",
X"05",
X"04",
X"04",
X"04",
X"03",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"02",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"05",
X"05",
X"05",
X"04",
X"05",
X"04",
X"05",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"01",
X"06",
X"04",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"04",
X"05",
X"05",
X"04",
X"05",
X"04",
X"05",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"06",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"04",
X"05",
X"05",
X"05",
X"05",
X"04",
X"05",
X"02",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"03",
X"05",
X"04",
X"05",
X"04",
X"04",
X"04",
X"03",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"02",
X"05",
X"04",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"05",
X"05",
X"05",
X"04",
X"05",
X"04",
X"05",
X"01",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"01",
X"06",
X"04",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"04",
X"05",
X"05",
X"04",
X"05",
X"04",
X"05",
X"02",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"06",
X"04",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"05",
X"05",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"01",
X"05",
X"04",
X"05",
X"04",
X"04",
X"05",
X"02",
X"FD",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"04",
X"05",
X"05",
X"04",
X"05",
X"04",
X"05",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"05",
X"04",
X"05",
X"04",
X"04",
X"05",
X"03",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"03",
X"05",
X"05",
X"05",
X"05",
X"04",
X"05",
X"00",
X"FD",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FE",
X"00",
X"05",
X"05",
X"05",
X"04",
X"05",
X"04",
X"04",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"FE",
X"00",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"01",
X"03",
X"02",
X"03",
X"02",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"02",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"03",
X"01",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"02",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"01",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"02",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"03",
X"03",
X"02",
X"03",
X"02",
X"03",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"03",
X"01",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"02",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"02",
X"03",
X"02",
X"02",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"01",
X"03",
X"02",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"02",
X"03",
X"03",
X"02",
X"03",
X"02",
X"02",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"01",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"01",
X"03",
X"02",
X"03",
X"02",
X"03",
X"02",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"02",
X"03",
X"02",
X"02",
X"02",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"00",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"

  );

  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;
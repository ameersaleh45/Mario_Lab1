--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bumb_sound is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(11 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end bumb_sound;

architecture arch of bumb_sound is

type table_type is array(0 to 4095) of std_logic_vector(7 downto 0);
signal sin_table : table_type;

begin

  SinTableTC_proc: process(RESET_N, CLK)
    constant sin_table : table_type := (

X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1D",
X"25",
X"22",
X"23",
X"21",
X"22",
X"20",
X"20",
X"1F",
X"1F",
X"1E",
X"1E",
X"1D",
X"1D",
X"1C",
X"1C",
X"1C",
X"1B",
X"1B",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"11",
X"10",
X"10",
X"0F",
X"10",
X"0E",
X"10",
X"0D",
X"11",
X"FB",
X"E8",
X"ED",
X"EA",
X"ED",
X"EB",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EF",
X"EE",
X"EF",
X"EF",
X"F0",
X"EF",
X"F0",
X"F0",
X"F1",
X"F0",
X"F1",
X"F1",
X"F2",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F5",
X"00",
X"1D",
X"19",
X"1B",
X"19",
X"1A",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"08",
X"EA",
X"E7",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F5",
X"F8",
X"F3",
X"06",
X"1D",
X"18",
X"1A",
X"18",
X"19",
X"17",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"16",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"08",
X"0B",
X"02",
X"E5",
X"E7",
X"E6",
X"E7",
X"E7",
X"E8",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F6",
X"14",
X"1B",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"09",
X"0A",
X"08",
X"0A",
X"07",
X"0C",
X"F4",
X"E2",
X"E7",
X"E5",
X"E7",
X"E6",
X"E8",
X"E7",
X"E9",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F4",
X"00",
X"1C",
X"18",
X"1A",
X"18",
X"19",
X"17",
X"18",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"15",
X"14",
X"14",
X"13",
X"13",
X"12",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"0A",
X"05",
X"E7",
X"E6",
X"E6",
X"E7",
X"E7",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F6",
X"14",
X"1C",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"07",
X"0A",
X"F1",
X"E2",
X"E6",
X"E4",
X"E7",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F9",
X"F4",
X"08",
X"1E",
X"18",
X"1B",
X"18",
X"1A",
X"18",
X"18",
X"17",
X"18",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"07",
X"0B",
X"FD",
X"E2",
X"E6",
X"E4",
X"E7",
X"E5",
X"E7",
X"E6",
X"E8",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F8",
X"F5",
X"FE",
X"1B",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"07",
X"08",
X"07",
X"08",
X"06",
X"0A",
X"FC",
X"E1",
X"E5",
X"E3",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F5",
X"02",
X"1E",
X"1A",
X"1C",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"08",
X"06",
X"09",
X"FF",
X"E2",
X"E5",
X"E4",
X"E5",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F6",
X"00",
X"1D",
X"1A",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"08",
X"06",
X"09",
X"00",
X"E3",
X"E5",
X"E4",
X"E5",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"00",
X"1E",
X"1B",
X"1C",
X"1B",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"07",
X"05",
X"08",
X"00",
X"E2",
X"E4",
X"E3",
X"E4",
X"E4",
X"E5",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E7",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"00",
X"1D",
X"1B",
X"1C",
X"1B",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"07",
X"07",
X"06",
X"07",
X"06",
X"07",
X"05",
X"08",
X"00",
X"E2",
X"E4",
X"E3",
X"E4",
X"E4",
X"E5",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E7",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F7",
X"F6",
X"F8",
X"F6",
X"F9",
X"F4",
X"0A",
X"1E",
X"19",
X"1B",
X"19",
X"1A",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"15",
X"16",
X"15",
X"15",
X"14",
X"14",
X"13",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"07",
X"EA",
X"E2",
X"E5",
X"E4",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F6",
X"00",
X"1D",
X"1A",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"09",
X"08",
X"08",
X"07",
X"08",
X"07",
X"09",
X"06",
X"0A",
X"F4",
X"E1",
X"E6",
X"E3",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"16",
X"1C",
X"1A",
X"1B",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"08",
X"08",
X"07",
X"08",
X"07",
X"08",
X"06",
X"09",
X"00",
X"E2",
X"E5",
X"E4",
X"E5",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F6",
X"F9",
X"F5",
X"0B",
X"1E",
X"19",
X"1C",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"07",
X"08",
X"07",
X"06",
X"E9",
X"E3",
X"E5",
X"E4",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F7",
X"F9",
X"F6",
X"00",
X"1D",
X"1A",
X"1B",
X"1A",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"17",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"06",
X"E8",
X"E4",
X"E6",
X"E6",
X"E6",
X"E7",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F6",
X"F8",
X"F5",
X"FE",
X"1B",
X"19",
X"1A",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"0A",
X"08",
X"0A",
X"08",
X"0A",
X"07",
X"0B",
X"FC",
X"E2",
X"E7",
X"E4",
X"E7",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F5",
X"F7",
X"F5",
X"F8",
X"F4",
X"0A",
X"1D",
X"18",
X"1B",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"08",
X"09",
X"07",
X"0A",
X"EE",
X"E3",
X"E7",
X"E5",
X"E7",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EC",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F9",
X"17",
X"1B",
X"19",
X"19",
X"19",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"16",
X"15",
X"15",
X"15",
X"14",
X"14",
X"14",
X"13",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"09",
X"08",
X"09",
X"07",
X"0A",
X"01",
X"E4",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F5",
X"F7",
X"F5",
X"F7",
X"F5",
X"F8",
X"F4",
X"03",
X"1D",
X"18",
X"1A",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"0A",
X"09",
X"0A",
X"08",
X"0A",
X"08",
X"0A",
X"07",
X"0B",
X"F5",
X"E2",
X"E7",
X"E4",
X"E7",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E8",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F8",
X"F5",
X"11",
X"1C",
X"18",
X"1A",
X"18",
X"19",
X"18",
X"18",
X"17",
X"17",
X"16",
X"16",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0F",
X"0F",
X"0E",
X"0E",
X"0E",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0B",
X"0B",
X"0B",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"0A",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"08",
X"08",
X"07",
X"E9",
X"E4",
X"E6",
X"E5",
X"E6",
X"E6",
X"E7",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"12",
X"1B",
X"17",
X"19",
X"17",
X"18",
X"16",
X"17",
X"16",
X"16",
X"15",
X"15",
X"14",
X"14",
X"14",
X"14",
X"13",
X"13",
X"12",
X"12",
X"12",
X"12",
X"11",
X"11",
X"11",
X"11",
X"10",
X"10",
X"10",
X"10",
X"0F",
X"0F",
X"0E",
X"0F",
X"0E",
X"0E",
X"0D",
X"0E",
X"0D",
X"0D",
X"0D",
X"0D",
X"0C",
X"0C",
X"0C",
X"0C",
X"0B",
X"0C",
X"0B",
X"0B",
X"0A",
X"0B",
X"0A",
X"0B",
X"09",
X"0A",
X"09",
X"0A",
X"08",
X"0B",
X"F1",
X"E3",
X"E8",
X"E6",
X"E8",
X"E7",
X"E8",
X"E8",
X"E9",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EB",
X"EB",
X"EB",
X"EB",
X"EC",
X"EC",
X"ED",
X"ED",
X"ED",
X"ED",
X"EE",
X"EE",
X"EE",
X"EF",
X"EF",
X"EF",
X"F0",
X"F0",
X"F0",
X"F0",
X"F1",
X"F1",
X"F1",
X"F1",
X"F2",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F5",
X"F5",
X"F5",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00"

);

  begin

    if (RESET_N='0') then
      Q <= sin_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sin_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;